`timescale 1ns / 1ps
module encoder(
    
    );
endmodule
